.title KiCad schematic
U3 Net-_C5-Pad1_ /TX /RX /2_INT0_ /3_INT1_ /_PD4_ +5V GND /XTAL1 /XTAL2 /5_PD5_ /_PD6_ /_PD7_ NC_01 /9_CE_ /10_CS_ /MOSI /MISO /SCK +5V NC_02 GND NC_03 NC_04 NC_05 NC_06 /SDA /SCL ATmega328-PU
C4 /XTAL1 GND 22p
C2 /XTAL2 GND 22p
C8 +5V GND 47uF
J2 /MISO +5V /SCK /MOSI Net-_C5-Pad1_ GND AVR-ISP-6
R2 +5V Net-_C5-Pad1_ 10k
R1 /XTAL1 /XTAL2 1M
D1 +5V Net-_C5-Pad1_ 1N4145
C9 +5V GND 100n
U1 GND +3V3 /9_CE_ /10_CS_ /SCK /MOSI /MISO /2_INT0_ NRF24L01_Breakout
J1 NEUT Net-_F1-Pad2_ 220V
U2 +3V3 GND +5V L78L33_TO92
C3 +5V GND 100n
C7 +3V3 GND 100n
C6 +3V3 GND 47uF
K1 LINE +5V Net-_J6-Pad1_ NC_07 Net-_D2-Pad2_ SANYOU_SRD_Form_C
D2 +5V Net-_D2-Pad2_ 1N4007
Q1 Net-_D2-Pad2_ Net-_Q1-Pad2_ GND BC547
R6 Net-_D6-Pad1_ Net-_Q1-Pad2_ 10k
D6 Net-_D6-Pad1_ /5_PD5_ 1N4148
J6 Net-_J6-Pad1_ NEUT LAMP
J3 +5V /3_INT1_ GND PIR
J4 +3V3 GND /SCL /SDA NC_08 BH1750
C1 +5V GND 220uF
F1 LINE Net-_F1-Pad2_ 500mA
Y1 /XTAL2 /XTAL1 Crystal
D3 Net-_D3-Pad1_ +5V red
D4 Net-_D4-Pad1_ +5V green
D5 Net-_D5-Pad1_ +5V yellow
R3 Net-_D3-Pad1_ /_PD4_ 470
R4 Net-_D4-Pad1_ /_PD6_ 470
R5 Net-_D5-Pad1_ /_PD7_ 470
SW1 GND Net-_C5-Pad1_ SW_Push
PS1 LINE NEUT GND +5V HLK-PM01
PS2 LINE NEUT +5V GND AC_DC_5V_3W-Converter_ACDC
H1 GND H
H2 GND H
H3 GND H
H4 MountingHole
J5 GND GND +5V /TX /RX /DTR FTDI
C5 Net-_C5-Pad1_ /DTR 100n
.end
